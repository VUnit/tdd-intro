package string_pkg is
   function to_string (data : integer_vector) return string;
end package;

package body string_pkg is
   function to_string (data : integer_vector) return string is
   begin
    return "";
  end function;
end package body;
