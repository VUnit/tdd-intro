package incrementer_pkg is
  constant increment_reg_addr : natural := 0;
end package incrementer_pkg;
